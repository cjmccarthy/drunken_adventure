--
-- VHDL Architecture ece411.SEXT5.untitled
--
-- Created:
--          by - mccart18.ews (gelib-057-16.ews.illinois.edu)
--          at - 03:45:36 03/12/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY SEXT5 IS
   PORT( 
      IR5down      : IN     LC3B_IMM5;
      offset5_SEXT : OUT    LC3B_WORD
   );

-- Declarations

END SEXT5 ;

--
ARCHITECTURE untitled OF SEXT5 IS
BEGIN
  offset5_SEXT <= IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down(4) & IR5down after DELAY_MUX2;
END ARCHITECTURE untitled;

