--
-- VHDL Architecture ece411.REG32.untitled
--
-- Created:
--          by - mccart18.ews (evrt-252-12.ews.illinois.edu)
--          at - 20:14:21 03/14/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY REG32 IS
-- Declarations

END REG32 ;

--
ARCHITECTURE untitled OF REG32 IS
BEGIN
END ARCHITECTURE untitled;

