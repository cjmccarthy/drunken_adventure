--
-- VHDL Architecture ece411.OWordJoinerH.untitled
--
-- Created:
--          by - hyunyi1.ews (evrt-252-10.ews.illinois.edu)
--          at - 20:46:18 03/27/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY OWordJoinerH IS
   PORT( 
      OWordIn   : IN     lc3b_oword;
      WordOut7  : IN     LC3B_WORD;
      OWordHOut : OUT    lc3b_oword
   );

-- Declarations

END OWordJoinerH ;

--
ARCHITECTURE untitled OF OWordJoinerH IS
BEGIN
  PROCESS(OWORDIN, WORDOUT7)
  variable TEMPOWORD :lc3b_oword;
  BEGIN
  tempoword:=OWORDIN;
  tempoword(127 downto 112):=wordout7;
  owordHout<=tempoword;
END PROCESS;
END ARCHITECTURE untitled;

