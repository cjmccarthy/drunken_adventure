--
-- VHDL Architecture ece411.OWordJoinerA.untitled
--
-- Created:
--          by - hyunyi1.ews (evrt-252-10.ews.illinois.edu)
--          at - 20:32:52 03/27/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY OWordJoinerA IS
   PORT( 
      OWordIn  : IN     lc3b_oword;
      WordOut  : IN     LC3B_WORD;
      OWordAOut: OUT    lc3b_oword
   );

-- Declarations

END OWORDJOINERA ;

--
ARCHITECTURE untitled OF OWORDJOINERA IS
BEGIN
  PROCESS(OWORDIN, WORDOUT)
  variable TEMPOWORD :lc3b_oword;
  BEGIN
  tempoword:=OWORDIN;
  tempoword(15 downto 0):=wordout;
  owordAout<=tempoword;
END PROCESS;
END ARCHITECTURE untitled;
